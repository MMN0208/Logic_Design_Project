module Part2 (SW, KEY, LEDR, HEX0, HEX2, HEX4, HEX5);
	input [8:0] SW;
	output [1:0] KEY;
	
	
endmodule