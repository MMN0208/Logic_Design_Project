module part1 (CLOCK_50, SW, KEY, LEDR, HEX0);
	input CLOCK_50;
	input [9:0] SW;
	input [1:0] KEY;
	output [9:0] LEDR;
	output [6:0] HEX0;
	
	
endmodule